`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module: Half_Adder
//////////////////////////////////////////////////////////////////////////////////

module Half_Adder(
    input A,
    input B,
    output Sum,
    output Cout
    );
    
    xor x1(Sum,A,B);
    and a1(Cout,A,B);
    
endmodule
